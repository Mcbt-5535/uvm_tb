class s12 extends s1#(abvasda);
sad wire 
213 1
d adsf 

 dasf;