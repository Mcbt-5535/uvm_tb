class t2 extends base_t;
dasf 231
123
dsf areg
123123 
