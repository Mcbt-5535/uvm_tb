class v22 extends v2;
typedef struct packed {
    
} 
231
3
sdas
;