class t123 extends t12;
sadasd
12312
dsf
import React from 'react'