class v21 extends v22;
adsf

fgdh
23
fds
