class v2 extends base_v;
adsf aa

adf 
 dasfasdfa dasfasdf

 dasfasdf
 fd 
