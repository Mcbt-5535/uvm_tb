class base_s extends uvm_sequence#(test1);
asda dasf
asda while () begin
    
    ``12`
    `4
end