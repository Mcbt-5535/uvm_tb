class base_v extends uvm_sequence;

dsa

dsada
asd

asd instance_name (.*);