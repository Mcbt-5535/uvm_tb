class base_t extends uvm_test;
adsf a

431325
32
423 
import React from 'react'