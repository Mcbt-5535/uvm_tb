class s2 extends base_s;
asdf asd
 3re
  1324

   fddg always_ff @( 
    
    ) begin : blockName
    
   end