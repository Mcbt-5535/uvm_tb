class t12 extends t1;
dsa dasf
213123

sada dasfasdf
1231