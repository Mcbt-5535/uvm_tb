class t1 extends uvm_test;
312
sewr;
sadasd

2313
import React from 'react'