class s1 extends uvm_sequence;
sadad aa
import React from 'react'

endclass