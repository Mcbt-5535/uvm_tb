class v1 extends uvm_sequence;
dasfasdf 
fgdh
 asd
 fgdha 
 ce_name (.*);