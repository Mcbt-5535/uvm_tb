class s123 extends s12#(123312,213123);
qewr qwer qsfdaSD
import React from 'react';
SAD qweqw 